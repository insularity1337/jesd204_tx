module rx_env (
  input               QPLL_REFCLK,
  input               DRPCLK     ,
  input               ACLK       ,
  input               ARESETN    ,
  input  [11:0]       AWADDR     ,
  input               AWVALID    ,
  output              AWREADY    ,
  input  [31:0]       WDATA      ,
  input  [ 3:0]       WSTRB      ,
  input               WVALID     ,
  output              WREADY     ,
  output [ 1:0]       BRESP      ,
  output              BVALID     ,
  input               BREADY     ,
  input  [11:0]       ARADDR     ,
  input               ARVALID    ,
  output              ARREADY    ,
  output [31:0]       RDATA      ,
  output [ 1:0]       RRESP      ,
  output              RVALID     ,
  input               RREADY     ,
  input               SYS_RESET  ,
  input               CLK        ,
  input               RST        ,
  input               SYSREF     ,
  output              SYNC_n     ,
  output              RX_ARESETN ,
  output              RX_TVALID  ,
  output [ 3:0][31:0] RX_TDATA   ,
  input  [ 3:0]       RX_N       ,
  input  [ 3:0]       RX_P
);

  logic rx_core_clk;

  logic [3:0][63:0] gt_rxdata      ;
  logic [3:0][ 3:0] gt_rxcharisk   ;
  logic [3:0][ 3:0] gt_rxdisperr   ;
  logic [3:0][ 3:0] gt_rxnotintable;
  logic [3:0][ 1:0] gt_rxheader    ;
  logic [3:0]       gt_rxmisalign  ;
  logic [3:0]       gt_rxblock_sync;

  jesd204b_rx link (
    .s_axi_aclk      (ACLK              ),
    .s_axi_aresetn   (ARESETN           ),
    .s_axi_awaddr    (AWADDR            ),
    .s_axi_awvalid   (AWVALID           ),
    .s_axi_awready   (AWREADY           ),
    .s_axi_wdata     (WDATA             ),
    .s_axi_wstrb     (WSTRB             ),
    .s_axi_wvalid    (WVALID            ),
    .s_axi_wready    (WREADY            ),
    .s_axi_bresp     (BRESP             ),
    .s_axi_bvalid    (BVALID            ),
    .s_axi_bready    (BREADY            ),
    .s_axi_araddr    (ARADDR            ),
    .s_axi_arvalid   (ARVALID           ),
    .s_axi_arready   (ARREADY           ),
    .s_axi_rdata     (RDATA             ),
    .s_axi_rresp     (RRESP             ),
    .s_axi_rvalid    (RVALID            ),
    .s_axi_rready    (RREADY            ),
    .rx_core_clk     (QPLL_REFCLK       ),
    .rx_core_reset   (RST               ),
    .rx_sysref       (SYSREF            ),
    .irq             (                  ),
    .rx_tdata        (RX_TDATA          ),
    .rx_tvalid       (RX_TVALID         ),
    .rx_aresetn      (RX_ARESETN        ),
    .rx_sof          (                  ),
    .rx_somf         (                  ),
    .rx_frm_err      (                  ),
    .rx_sync         (SYNC_n            ),
    .encommaalign    (rxencommaalign    ),
    .rx_reset_gt     (rx_reset_gt       ),
    .rx_reset_done   (rx_reset_done     ),
    .gt0_rxdata      (gt_rxdata[0]      ),
    .gt0_rxcharisk   (gt_rxcharisk[0]   ),
    .gt0_rxdisperr   (gt_rxdisperr[0]   ),
    .gt0_rxnotintable(gt_rxnotintable[0]),
    .gt0_rxheader    (gt_rxheader[0]    ),
    .gt0_rxmisalign  (gt_rxmisalign[0]  ),
    .gt0_rxblock_sync(gt_rxblock_sync[0]),
    .gt1_rxdata      (gt_rxdata[1]      ),
    .gt1_rxcharisk   (gt_rxcharisk[1]   ),
    .gt1_rxdisperr   (gt_rxdisperr[1]   ),
    .gt1_rxnotintable(gt_rxnotintable[1]),
    .gt1_rxheader    (gt_rxheader[1]    ),
    .gt1_rxmisalign  (gt_rxmisalign[1]  ),
    .gt1_rxblock_sync(gt_rxblock_sync[1]),
    .gt2_rxdata      (gt_rxdata[2]      ),
    .gt2_rxcharisk   (gt_rxcharisk[2]   ),
    .gt2_rxdisperr   (gt_rxdisperr[2]   ),
    .gt2_rxnotintable(gt_rxnotintable[2]),
    .gt2_rxheader    (gt_rxheader[2]    ),
    .gt2_rxmisalign  (gt_rxmisalign[2]  ),
    .gt2_rxblock_sync(gt_rxblock_sync[2]),
    .gt3_rxdata      (gt_rxdata[3]      ),
    .gt3_rxcharisk   (gt_rxcharisk[3]   ),
    .gt3_rxdisperr   (gt_rxdisperr[3]   ),
    .gt3_rxnotintable(gt_rxnotintable[3]),
    .gt3_rxheader    (gt_rxheader[3]    ),
    .gt3_rxmisalign  (gt_rxmisalign[3]  ),
    .gt3_rxblock_sync(gt_rxblock_sync[3])
  );

  jesd204b_rx_phy phy (
    .qpll0_refclk            (QPLL_REFCLK       ),
    .drpclk                  (DRPCLK            ),
    .tx_reset_gt             (rx_reset_gt       ),
    .rx_reset_gt             (rx_reset_gt       ),
    .tx_sys_reset            (SYS_RESET         ),
    .rx_sys_reset            (SYS_RESET         ),
    .txp_out                 (                  ),
    .txn_out                 (                  ),
    .rxp_in                  (RX_P              ),
    .rxn_in                  (RX_N              ),
    .tx_core_clk             (QPLL_REFCLK       ),
    .rx_core_clk             (QPLL_REFCLK       ),
    .txoutclk                (txoutclk          ),
    .rxoutclk                (rxoutclk          ),
    .gt_prbssel              (4'h0              ),
    .gt0_txdata              (32'h00000000      ),
    .gt0_txcharisk           (4'h0              ),
    .tx_reset_done           (tx_reset_done     ),
    .gt_powergood            (gt_powergood      ),
    .gt0_rxdata              (gt_rxdata[0]      ),
    .gt0_rxcharisk           (gt_rxcharisk[0]   ),
    .gt0_rxdisperr           (gt_rxdisperr[0]   ),
    .gt0_rxnotintable        (gt_rxnotintable[0]),
    .gt1_rxdata              (gt_rxdata[1]      ),
    .gt1_rxcharisk           (gt_rxcharisk[1]   ),
    .gt1_rxdisperr           (gt_rxdisperr[1]   ),
    .gt1_rxnotintable        (gt_rxnotintable[1]),
    .gt2_rxdata              (gt_rxdata[2]      ),
    .gt2_rxcharisk           (gt_rxcharisk[2]   ),
    .gt2_rxdisperr           (gt_rxdisperr[2]   ),
    .gt2_rxnotintable        (gt_rxnotintable[2]),
    .gt3_rxdata              (gt_rxdata[3]      ),
    .gt3_rxcharisk           (gt_rxcharisk[3]   ),
    .gt3_rxdisperr           (gt_rxdisperr[3]   ),
    .gt3_rxnotintable        (gt_rxnotintable[3]),
    .rx_reset_done           (rx_reset_done     ),
    .rxencommaalign          (rxencommaalign    ),
    .common0_qpll0_clk_out   (                  ),
    .common0_qpll0_refclk_out(                  ),
    .common0_qpll0_lock_out  (                  )
  );

endmodule